////////////////////////////////////////////////////////////////////////////////
//                                            __ _      _     _               //
//                                           / _(_)    | |   | |              //
//                __ _ _   _  ___  ___ _ __ | |_ _  ___| | __| |              //
//               / _` | | | |/ _ \/ _ \ '_ \|  _| |/ _ \ |/ _` |              //
//              | (_| | |_| |  __/  __/ | | | | | |  __/ | (_| |              //
//               \__, |\__,_|\___|\___|_| |_|_| |_|\___|_|\__,_|              //
//                  | |                                                       //
//                  |_|                                                       //
//                                                                            //
//                                                                            //
//              MSP430 CPU                                                    //
//              Processing Unit                                               //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

/* Copyright (c) 2015-2016 by the author(s)
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 *
 * =============================================================================
 * Author(s):
 *   Francisco Javier Reina Campo <frareicam@gmail.com>
 */

module  msp430_template08 (
  // OUTPUTs
  output      [15:0] per_dout,        // Peripheral data output

  // INPUTs
  input              mclk,            // Main system clock
  input       [13:0] per_addr,        // Peripheral address
  input       [15:0] per_din,         // Peripheral data input
  input              per_en,          // Peripheral enable (high active)
  input        [1:0] per_we,          // Peripheral write enable (high active)
  input              puc_rst          // Main system reset
);

  //=============================================================================
  // 1)  PARAMETER DECLARATION
  //=============================================================================

  // Register base address (must be aligned to decoder bit width)
  parameter       [14:0] BASE_ADDR   = 15'h0090;

  // Decoder bit width (defines how many bits are considered for address decoding)
  parameter              DEC_WD      =  2;

  // Register addresses offset
  parameter [DEC_WD-1:0] CNTRL1      =  'h0,
  CNTRL2      =  'h1,
  CNTRL3      =  'h2,
  CNTRL4      =  'h3;

  // Register one-hot decoder utilities
  parameter              DEC_SZ      =  (1 << DEC_WD);
  parameter [DEC_SZ-1:0] BASE_REG    =  {{DEC_SZ-1{1'b0}}, 1'b1};

  // Register one-hot decoder
  parameter [DEC_SZ-1:0] CNTRL1_D  = (BASE_REG << CNTRL1),
  CNTRL2_D  = (BASE_REG << CNTRL2), 
  CNTRL3_D  = (BASE_REG << CNTRL3), 
  CNTRL4_D  = (BASE_REG << CNTRL4); 

  //============================================================================
  // 2)  REGISTER DECODER
  //============================================================================

  // Local register selection
  wire              reg_sel      =  per_en & (per_addr[13:DEC_WD-1]==BASE_ADDR[14:DEC_WD]);

  // Register local address
  wire [DEC_WD-1:0] reg_addr     =  {1'b0, per_addr[DEC_WD-2:0]};

  // Register address decode
  wire [DEC_SZ-1:0] reg_dec      = (CNTRL1_D  &  {DEC_SZ{(reg_addr==(CNTRL1 >>1))}}) |
                                   (CNTRL2_D  &  {DEC_SZ{(reg_addr==(CNTRL2 >>1))}}) |
                                   (CNTRL3_D  &  {DEC_SZ{(reg_addr==(CNTRL3 >>1))}}) |
                                   (CNTRL4_D  &  {DEC_SZ{(reg_addr==(CNTRL4 >>1))}});

  // Read/Write probes
  wire              reg_lo_write =  per_we[0] & reg_sel;
  wire              reg_hi_write =  per_we[1] & reg_sel;
  wire              reg_read     = ~|per_we   & reg_sel;

  // Read/Write vectors
  wire [DEC_SZ-1:0] reg_hi_wr    = reg_dec & {DEC_SZ{reg_hi_write}};
  wire [DEC_SZ-1:0] reg_lo_wr    = reg_dec & {DEC_SZ{reg_lo_write}};
  wire [DEC_SZ-1:0] reg_rd       = reg_dec & {DEC_SZ{reg_read}};

  //============================================================================
  // 3) REGISTERS
  //============================================================================

  // CNTRL1 Register
  //-----------------
  reg  [7:0] cntrl1;

  wire       cntrl1_wr  = CNTRL1[0] ? reg_hi_wr[CNTRL1] : reg_lo_wr[CNTRL1];
  wire [7:0] cntrl1_nxt = CNTRL1[0] ? per_din[15:8]     : per_din[7:0];

  always @ (posedge mclk or posedge puc_rst) begin
    if (puc_rst)        cntrl1 <=  8'h00;
    else if (cntrl1_wr) cntrl1 <=  cntrl1_nxt;
  end

  // CNTRL2 Register
  //-----------------
  reg  [7:0] cntrl2;

  wire       cntrl2_wr  = CNTRL2[0] ? reg_hi_wr[CNTRL2] : reg_lo_wr[CNTRL2];
  wire [7:0] cntrl2_nxt = CNTRL2[0] ? per_din[15:8]     : per_din[7:0];

  always @ (posedge mclk or posedge puc_rst) begin
    if (puc_rst)        cntrl2 <=  8'h00;
    else if (cntrl2_wr) cntrl2 <=  cntrl2_nxt;
  end

  // CNTRL3 Register
  //-----------------
  reg  [7:0] cntrl3;

  wire       cntrl3_wr  = CNTRL3[0] ? reg_hi_wr[CNTRL3] : reg_lo_wr[CNTRL3];
  wire [7:0] cntrl3_nxt = CNTRL3[0] ? per_din[15:8]     : per_din[7:0];

  always @ (posedge mclk or posedge puc_rst) begin
    if (puc_rst)        cntrl3 <=  8'h00;
    else if (cntrl3_wr) cntrl3 <=  cntrl3_nxt;
  end

  // CNTRL4 Register
  //-----------------
  reg  [7:0] cntrl4;

  wire       cntrl4_wr  = CNTRL4[0] ? reg_hi_wr[CNTRL4] : reg_lo_wr[CNTRL4];
  wire [7:0] cntrl4_nxt = CNTRL4[0] ? per_din[15:8]     : per_din[7:0];

  always @ (posedge mclk or posedge puc_rst) begin
    if (puc_rst)        cntrl4 <=  8'h00;
    else if (cntrl4_wr) cntrl4 <=  cntrl4_nxt;
  end

  //============================================================================
  // 4) DATA OUTPUT GENERATION
  //============================================================================

  // Data output mux
  wire [15:0] cntrl1_rd   = {8'h00, (cntrl1  & {8{reg_rd[CNTRL1]}})}  << (8 & {4{CNTRL1[0]}});
  wire [15:0] cntrl2_rd   = {8'h00, (cntrl2  & {8{reg_rd[CNTRL2]}})}  << (8 & {4{CNTRL2[0]}});
  wire [15:0] cntrl3_rd   = {8'h00, (cntrl3  & {8{reg_rd[CNTRL3]}})}  << (8 & {4{CNTRL3[0]}});
  wire [15:0] cntrl4_rd   = {8'h00, (cntrl4  & {8{reg_rd[CNTRL4]}})}  << (8 & {4{CNTRL4[0]}});

  assign      per_dout  =  cntrl1_rd  |
                           cntrl2_rd  |
                           cntrl3_rd  |
                           cntrl4_rd;   
endmodule // msp430_template08
