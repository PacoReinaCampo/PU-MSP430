../../../../bench/verilog/baremetal/regression/leds.sv