../../../../../../../bench/verilog/baremetal/cases/leds.sv