../../../bench/verilog/regression/two-op_add.sv